// $Id: $
// File name:   bit_stuffer.sv
// Created:     2/26/2019
// Author:      Nur Nadhira Aqilah Binti Mohd Shah
// Lab Section: 2
// Version:     1.0  Initial Design Entry
// Description: bit stuffer for usb tx

module tx_bit_stuffer
(
    input wire clk,
    input wire n_rst,
    input wire shift_enable,
    input wire serial_out,
    output reg pause
    //output wire val
);
    //reg [15:0] prev_pause;
    wire count_enable;
    assign count_enable = serial_out & shift_enable;
    
    flex_counter #(
    	.NUM_CNT_BITS(3)
    )
    CORE (
	.clk(clk),
	.n_rst(n_rst),
	.clear(!serial_out),
	.count_enable(count_enable),
	.rollover_val(3'd5),
	.count_out(),
	.rollover_flag(pause)
    );
    
 /*   always_ff @ (posedge clk, negedge n_rst) begin
        if (!n_rst) begin
        	prev_pause <= 1'b0;
        end
	else begin
        	prev_pause[0] <= prev_pause[1];
        	prev_pause[1] <= prev_pause[2];
        	prev_pause[2] <= prev_pause[3];
        	prev_pause[3] <= prev_pause[4];
        	prev_pause[4] <= prev_pause[5];
        	prev_pause[5] <= prev_pause[6];
        	prev_pause[6] <= prev_pause[7];
        	prev_pause[7] <= prev_pause[8];
        	prev_pause[8] <= prev_pause[9];
        	prev_pause[9] <= prev_pause[10];
        	prev_pause[10] <= prev_pause[11];
        	prev_pause[11] <= prev_pause[12];
        	prev_pause[12] <= prev_pause[13];
        	prev_pause[13] <= prev_pause[14];
        	prev_pause[14] <= prev_pause[15];
	        prev_pause[15] <= pause;
        end
    end
    assign val = prev_pause[15];
*/


endmodule

